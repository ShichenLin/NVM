package nvm_pkg();

endpackage
