`include "gc_controller_if.vh"

module gc_controller(
	gc_controller_if.gcc gccif
);

endmodule
