`include "garbage_collection_if.vh"

module garbage_collection(
	input logic CLK, nRST,
	garbage_collection_if.gc gcif
);


endmodule
